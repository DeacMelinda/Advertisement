library ieee;
use ieee.std_logic_1164.all;

entity copiere is
	port(A1, A2, A3, A4: in std_logic_vector(6 downto 0);
	C1, C2, C3, C4, en: in std_logic;
	B: out std_logic_vector(6 downto 0));
end copiere;



architecture copiere of copiere is	   
signal aux: std_logic_vector(6 downto 0);
begin
	
			
end copiere;


